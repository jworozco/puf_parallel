package puf_pkg;
    typedef enum logic [1:0] { START, PUF1, PUF2, HALT } state_t;
endpackage
